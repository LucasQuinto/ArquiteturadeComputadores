<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>3,9,132.8,-64.7</PageViewport>
<gate>
<ID>2</ID>
<type>AA_TOGGLE</type>
<position>7,-5.5</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>15,-7.5</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>7,-11.5</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_TOGGLE</type>
<position>14.5,-13</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_AND2</type>
<position>35.5,-7</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_AND2</type>
<position>35.5,-18</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>7 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_AND2</type>
<position>35.5,-28.5</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_AND2</type>
<position>55.5,-33.5</position>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>8 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>24</ID>
<type>AA_AND2</type>
<position>41.5,-49</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>7 </input>
<output>
<ID>OUT</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>28</ID>
<type>GA_LED</type>
<position>98.5,-5</position>
<input>
<ID>N_in2</ID>17 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>30</ID>
<type>GA_LED</type>
<position>107,-5</position>
<input>
<ID>N_in2</ID>15 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>32</ID>
<type>GA_LED</type>
<position>115,-5</position>
<input>
<ID>N_in2</ID>16 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>34</ID>
<type>GA_LED</type>
<position>124.5,-6.5</position>
<input>
<ID>N_in2</ID>4 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>36</ID>
<type>AI_XOR2</type>
<position>58,-16.5</position>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>8 </input>
<output>
<ID>OUT</ID>16 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>38</ID>
<type>AI_XOR2</type>
<position>75.5,-31.5</position>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_1</ID>11 </input>
<output>
<ID>OUT</ID>15 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>40</ID>
<type>AA_AND2</type>
<position>74,-50.5</position>
<input>
<ID>IN_0</ID>11 </input>
<input>
<ID>IN_1</ID>10 </input>
<output>
<ID>OUT</ID>17 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>42</ID>
<type>AA_LABEL</type>
<position>16.5,-4</position>
<gparam>LABEL_TEXT a1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>44</ID>
<type>AA_LABEL</type>
<position>7.5,-2</position>
<gparam>LABEL_TEXT a2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>46</ID>
<type>AA_LABEL</type>
<position>15.5,-16.5</position>
<gparam>LABEL_TEXT b1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>48</ID>
<type>AA_LABEL</type>
<position>7.5,-15</position>
<gparam>LABEL_TEXT b2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>50</ID>
<type>AA_LABEL</type>
<position>124,-3</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>52</ID>
<type>AA_LABEL</type>
<position>115,-1.5</position>
<gparam>LABEL_TEXT 2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>54</ID>
<type>AA_LABEL</type>
<position>107,-1.5</position>
<gparam>LABEL_TEXT 4</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>56</ID>
<type>AA_LABEL</type>
<position>98.5,-1.5</position>
<gparam>LABEL_TEXT 8</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>17,-7.5,32.5,-7.5</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>29 3</intersection>
<intersection>32.5 5</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>29,-27.5,29,-7.5</points>
<intersection>-27.5 4</intersection>
<intersection>-7.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>29,-27.5,32.5,-27.5</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>29 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>32.5,-7.5,32.5,-6</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>-7.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-13,24.5,-8</points>
<intersection>-13 2</intersection>
<intersection>-8 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24.5,-8,32.5,-8</points>
<connection>
<GID>10</GID>
<name>IN_1</name></connection>
<intersection>24.5 0</intersection>
<intersection>32.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16.5,-13,24.5,-13</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>24.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>32.5,-17,32.5,-8</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>-8 1</intersection></vsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124.5,-7.5,124.5,-7</points>
<connection>
<GID>34</GID>
<name>N_in2</name></connection>
<intersection>-7 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38.5,-7,124.5,-7</points>
<connection>
<GID>10</GID>
<name>OUT</name></connection>
<intersection>124.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20.5,-31,20.5,-11.5</points>
<intersection>-31 1</intersection>
<intersection>-11.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20.5,-31,38.5,-31</points>
<intersection>20.5 0</intersection>
<intersection>32.5 4</intersection>
<intersection>38.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>9,-11.5,20.5,-11.5</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>20.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>38.5,-48,38.5,-31</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>-31 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>32.5,-31,32.5,-29.5</points>
<connection>
<GID>14</GID>
<name>IN_1</name></connection>
<intersection>-31 1</intersection></vsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23.5,-50,23.5,-5.5</points>
<intersection>-50 1</intersection>
<intersection>-19 3</intersection>
<intersection>-5.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23.5,-50,38.5,-50</points>
<connection>
<GID>24</GID>
<name>IN_1</name></connection>
<intersection>23.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>9,-5.5,23.5,-5.5</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>23.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>23.5,-19,32.5,-19</points>
<connection>
<GID>12</GID>
<name>IN_1</name></connection>
<intersection>23.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44.5,-34.5,44.5,-17.5</points>
<intersection>-34.5 3</intersection>
<intersection>-25.5 2</intersection>
<intersection>-17.5 6</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>41.5,-25.5,44.5,-25.5</points>
<intersection>41.5 4</intersection>
<intersection>44.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>44.5,-34.5,52.5,-34.5</points>
<connection>
<GID>16</GID>
<name>IN_1</name></connection>
<intersection>44.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>41.5,-28.5,41.5,-25.5</points>
<intersection>-28.5 5</intersection>
<intersection>-25.5 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>38.5,-28.5,41.5,-28.5</points>
<connection>
<GID>14</GID>
<name>OUT</name></connection>
<intersection>41.5 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>44.5,-17.5,55,-17.5</points>
<connection>
<GID>36</GID>
<name>IN_1</name></connection>
<intersection>44.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44.5,-20.5,44.5,-20</points>
<intersection>-20.5 2</intersection>
<intersection>-20 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44.5,-20,54,-20</points>
<intersection>44.5 0</intersection>
<intersection>52.5 3</intersection>
<intersection>54 5</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>38.5,-20.5,44.5,-20.5</points>
<intersection>38.5 4</intersection>
<intersection>44.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>52.5,-32.5,52.5,-20</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>-20 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>38.5,-20.5,38.5,-18</points>
<connection>
<GID>12</GID>
<name>OUT</name></connection>
<intersection>-20.5 2</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>54,-20,54,-15.5</points>
<intersection>-20 1</intersection>
<intersection>-15.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>54,-15.5,55,-15.5</points>
<connection>
<GID>36</GID>
<name>IN_0</name></connection>
<intersection>54 5</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,-51,57,-49</points>
<intersection>-51 3</intersection>
<intersection>-49 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>44.5,-49,57,-49</points>
<connection>
<GID>24</GID>
<name>OUT</name></connection>
<intersection>57 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>57,-51,71,-51</points>
<intersection>57 0</intersection>
<intersection>69 4</intersection>
<intersection>71 5</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>69,-51,69,-30.5</points>
<intersection>-51 3</intersection>
<intersection>-30.5 6</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>71,-51.5,71,-51</points>
<connection>
<GID>40</GID>
<name>IN_1</name></connection>
<intersection>-51 3</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>69,-30.5,72.5,-30.5</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<intersection>69 4</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64,-33.5,64,-32.5</points>
<intersection>-33.5 2</intersection>
<intersection>-32.5 5</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>58.5,-33.5,64,-33.5</points>
<connection>
<GID>16</GID>
<name>OUT</name></connection>
<intersection>64 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>64,-32.5,72.5,-32.5</points>
<connection>
<GID>38</GID>
<name>IN_1</name></connection>
<intersection>64 0</intersection>
<intersection>71 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>71,-49.5,71,-32.5</points>
<connection>
<GID>40</GID>
<name>IN_0</name></connection>
<intersection>-32.5 5</intersection></vsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107,-31.5,107,-6</points>
<connection>
<GID>30</GID>
<name>N_in2</name></connection>
<intersection>-31.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>78.5,-31.5,107,-31.5</points>
<connection>
<GID>38</GID>
<name>OUT</name></connection>
<intersection>107 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115,-16.5,115,-6</points>
<connection>
<GID>32</GID>
<name>N_in2</name></connection>
<intersection>-16.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>61,-16.5,115,-16.5</points>
<connection>
<GID>36</GID>
<name>OUT</name></connection>
<intersection>115 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>98.5,-50.5,98.5,-6</points>
<connection>
<GID>28</GID>
<name>N_in2</name></connection>
<intersection>-50.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77,-50.5,98.5,-50.5</points>
<connection>
<GID>40</GID>
<name>OUT</name></connection>
<intersection>98.5 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,129.8,-73.7</PageViewport></page 1>
<page 2>
<PageViewport>0,0,129.8,-73.7</PageViewport></page 2>
<page 3>
<PageViewport>0,0,129.8,-73.7</PageViewport></page 3>
<page 4>
<PageViewport>0,0,129.8,-73.7</PageViewport></page 4>
<page 5>
<PageViewport>0,0,129.8,-73.7</PageViewport></page 5>
<page 6>
<PageViewport>0,0,129.8,-73.7</PageViewport></page 6>
<page 7>
<PageViewport>0,0,129.8,-73.7</PageViewport></page 7>
<page 8>
<PageViewport>0,0,129.8,-73.7</PageViewport></page 8>
<page 9>
<PageViewport>0,0,129.8,-73.7</PageViewport></page 9></circuit>